module imem(input  [31:0] addr,
            output [31:0] data);

  reg  [31:0] RAM[255:0];

  integer i;
  initial
    begin
      for (i = 0; i < 255; i = i + 1) begin
        RAM[i] = 0;
      end
      //$readmemh("memfile.dat",RAM);
/*      RAM[0]  = 32'b001000_00000_00001_0000000000000001; // addi r1, r0, 1
      RAM[1]  = 32'b001000_00000_00010_0000000000001011; // addi r2, r0, 11
      RAM[2]  = 32'b001000_00000_00011_0000000000000111; // addi r3, r0, 7

      RAM[3]  = 32'b001000_00001_00001_0000000000000001; // addi r1, r1, 1
      RAM[4]  = 32'b000101_00010_00001_0000000000000011; // bne r1, r2, 2
      RAM[5]  = 32'b101011_00000_00011_0000000000000100; // sw r3
      RAM[6]  = 32'b100011_00000_00001_0000000000000100; // lw r1
      RAM[7]  = 32'b000010_00000_00000_0000000000000111; // jump 
*/    

/*
      // Simple send  
      RAM[0]  = 32'b001000_00000_00001_0000000001001000; // addi r1, r0, 1
      RAM[1]  = 32'b101011_11111_00001_0000000000000001; // set tx byte
      RAM[2]  = 32'b001000_00000_00001_0000000000000001; // addi r1, r0, 1
      RAM[3]  = 32'b101011_11111_00001_0000000000000000; // set transmit
      RAM[4]  = 32'b101011_11111_00000_0000000000000000; // unset transmit
      RAM[5]  = 32'b000000_00000_00000_0000000000000000;
      RAM[6]  = 32'b000000_00000_00000_0000000000000000;
      RAM[7]  = 32'b000010_00000_00000_0000000000000111; // jump 
*/

      // Fibonacci
      RAM[0]  = 32'b001000_00000_00001_0000000000000001; // addi r1, r0, 1

      RAM[1]  = 32'b000000_00000_00001_00010_00000100000; // add r2, r0, r1
      RAM[2]  = 32'b001000_00001_00000_0000000000000000; // addi r0, r1, 0
      RAM[3]  = 32'b001000_00010_00001_0000000000000000; // addi r1, r2, 0

      RAM[4]  = 32'b101011_11111_00001_0000000000000001; // set tx byte
      RAM[5]  = 32'b001000_10000_10001_0000000000000001; // addi r1, r0, 1
      RAM[6]  = 32'b101011_11111_10001_0000000000000000; // set transmit
      RAM[7]  = 32'b101011_11111_10000_0000000000000000; // unset transmit

      //loop while transmission is in progress
      RAM[8]  = 32'b100011_11111_10011_0000000000000000; // lw r1
      RAM[9]  = 32'b000000_10011_10001_10011_00000100100; // and
      RAM[10] = 32'b000101_10000_10011_0000000000001000; // bne r1, r2, 2
      
      RAM[13] = 32'b000010_00000_00000_0000000000000001; // jump 
/*      // Echo
      RAM[0]  = 32'b001000_00000_00010_0000000000001010; // r2 := 10
      RAM[1]  = 32'b001000_00000_00011_0000000000000000; // r3 := 0
      RAM[2]  = 32'b001000_10000_10001_0000000000000001; // r17 := 1
     
      //store received chars to buffer
      RAM[7]  = 32'b001000_10000_10100_0000000000000010; // addi r1, r0, 1
      
      RAM[8]  = 32'b100011_11111_10011_0000000000000000; // lw r1
      RAM[9]  = 32'b000000_10011_10100_10011_00000100100; // and
      RAM[10] = 32'b000101_10100_10011_0000000000001000; // bne r1, r2, 2
      RAM[11] = 32'b100011_11111_00001_0000000000000001; // lw r1
      RAM[12] = 32'b101011_11111_10000_0000000000000010; // clear recv reg
      RAM[13] = 32'b101011_00011_00001_0000000000000000; // mem[r3] := r1
      RAM[14] = 32'b001000_00011_00011_0000000000000001; // r3 := r3 + 1
      RAM[15] = 32'b000101_00010_00001_0000000000001000; // bne r1, r2
     
      RAM[0]  = 32'b001000_00000_00001_0000000001001000; // addi r1, r0, 1
      RAM[1]  = 32'b101011_00000_00001_0000000000000000; // mem[r3] := r1
      RAM[2]  = 32'b101011_00000_00001_0000000000000001; // mem[r3+1] := r1
      RAM[3]  = 32'b101011_00000_00001_0000000000000010; // mem[r3+2] := r1
      RAM[4]  = 32'b001000_00000_00001_0000000000001010; // addi r1, r0, 1
      RAM[5]  = 32'b101011_00000_00001_0000000000000011; // mem[r3+2] := r1
      RAM[6]  = 32'b001000_10000_10001_0000000000000001; // addi r1, r0, 1
      RAM[7]  = 32'b001000_00000_00010_0000000000001010; // r2 := 10

      //send from buffer
      RAM[16] = 32'b001000_00000_00011_0000000000000000; // r3 := 0

      RAM[17] = 32'b100011_00011_00001_0000000000000000; // r1 := mem[r3]
      RAM[18] = 32'b101011_11111_00001_0000000000000001; // mem[tx_byte] := r1
      RAM[20] = 32'b101011_11111_10001_0000000000000000; // set transmit
      RAM[25] = 32'b101011_11111_10000_0000000000000000; // unset transmit

      //loop while transmission is in progress
      RAM[32] = 32'b100011_11111_10011_0000000000000000; // lw r1
      RAM[33] = 32'b000000_10011_10001_10011_00000100100; // and
      RAM[34] = 32'b000101_10000_10011_0000000000010110; // bne r1, r2, 2

      RAM[35] = 32'b001000_00011_00011_0000000000000001; // r3 := r3 + 1
     
      RAM[36] = 32'b000101_00010_00001_0000000000010001; // bne r1, r2
      
      RAM[40] = 32'b000010_00000_00000_0000000000101000; // jump 
*/    end
  assign data = RAM[addr];
endmodule
